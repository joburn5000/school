module aliens_rom
(
	input 	[7:0] addr,
	output 	[7:0] data
);

	logic[7:0] addr_reg;

	parameter [0:48][7:0] ROM = {

		8'b01000010, //0   crab
		8'b00100100, //1     
		8'b01111110, //2  
		8'b11011011, //3 
		8'b11111111, //4
		8'b10111101, //5  
		8'b10100101, //6 
		8'b00100100, //7 
		
		8'b01000010, //8   
		8'b10100101, //9     
		8'b10111101, //10  
		8'b11011011, //11 
		8'b11111111, //12
		8'b01111110, //13 
		8'b00100100, //14
		8'b01000010, //15  
		
		8'b00011000, //16   squid
		8'b00111100, //17   
		8'b01111110, //18  
		8'b11011011, //19  
		8'b11111111, //20  
		8'b01011010, //21  
		8'b10000001, //22  
		8'b01000010, //23
		
		8'b00011000, //24    
		8'b00111100, //25    
		8'b01111110, //26  
		8'b11011011, //27 
		8'b11111111, //28  
		8'b00100100, //29  
		8'b01011010, //30  
		8'b10100101, //31
		
		8'b00011000, //32   octopus
		8'b01111110, //33  
		8'b11111111, //34 
		8'b11011011, //35 
		8'b11111111, //36 
		8'b01100110, //37  
		8'b11011011, //38 
		8'b01100110, //39 
		
		8'b00011000, //40   
		8'b01111110, //41  
		8'b11111111, //42 
		8'b11011011, //43 
		8'b11111111, //44 
		8'b00100100, //45  
		8'b01011010, //46 
		8'b10000001, //47 
		
	};

	assign data = ROM[addr];
	
endmodule 